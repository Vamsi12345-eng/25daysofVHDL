
--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   10:59:54 01/13/2024
-- Design Name:   half_add
-- Module Name:   half_add_test.vhd
-- Project Name:  day_001
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: half_add
--
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends 
-- that these types always be used for the top-level I/O of a design in order 
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.all;
USE ieee.numeric_std.ALL;


ENTITY half_add_test_vhd IS
END half_add_test_vhd;

ARCHITECTURE behavior OF half_add_test_vhd IS 

	-- Component Declaration for the Unit Under Test (UUT)
	COMPONENT half_add
	PORT(
		a : IN std_logic;
		b : IN std_logic;          
		sum : OUT std_logic;
		carry : OUT std_logic
		);
	END COMPONENT;

	--Inputs
	SIGNAL a :  std_logic := '0';
	SIGNAL b :  std_logic := '0';

	--Outputs
	SIGNAL sum :  std_logic;
	SIGNAL carry :  std_logic;

BEGIN

	-- Instantiate the Unit Under Test (UUT)
	uut: half_add PORT MAP(
		a => a,
		b => b,
		sum => sum,
		carry => carry
	);

	tb : PROCESS
	BEGIN

    a <= '0';
	 b <= '1';
	 
	 wait for 10ns;
	 
	     a <= '1';
	 b <= '1';
	 
	 wait for 10ns;
	 
	 	     a <= '0';
	 b <= '0';
	 
	 wait for 10ns;
	 
	 	     a <= '1';
	 b <= '0';
	 
    wait;
	 

	END PROCESS;

END;
